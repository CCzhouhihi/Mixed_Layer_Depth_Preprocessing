netcdf HYCOMnwp_mask {
dimensions:
	time = UNLIMITED ; // (0 currently)
	latitude = 186 ;
	longitude = 53 ;
variables:
	float LANDMASK(time, latitude, longitude) ;
		LANDMASK:long_name = "LANDMASK 1 represents should be masked" ;
	double latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degree_north" ;
		latitude:axis = "Y" ;
	double longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degree_east" ;
		longitude:modulo = "360 degrees" ;
		longitude:axis = "X" ;
	double time(time) ;
		time:units = "hours since 2000-01-01 00:00:00" ;
		time:time_origin = "2000-01-01 00:00:00" ;
		time:calendar = "gregorian" ;
		time:axis = "T" ;

// global attributes:
		:TITILE = "MASK in Northwest Pacific" ;
}
